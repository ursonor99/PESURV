module top1(
      input wire clk

    );
s_core_pipelined uuts_core();

endmodule