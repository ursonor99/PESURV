module top1(
      input wire clk;
      input wire ok
    );
s_core_pipelined uuts_core();

endmodule